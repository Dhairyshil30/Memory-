`include "memory.v"

`include "comm.sv"
`include "interface.sv"
`include "mem_txs.sv"
`include "mem_asserstion.sv"

`include "mem_gen.sv"
`include "mem_bfm.sv"
`include "mem_mon.sv"
`include "mem_cov.sv"
`include "mem_sbd.sv"


`include "agent.sv"
`include "mem_env.sv"

`include "top.sv"

